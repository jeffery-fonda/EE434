
.GLOBAL VDD
.GLOBAL VSS

.SUBCKT myInv_X1 A ZN VDD VSS
mn1 ZN A VSS VSS NMOS_HP L=0.05u W=0.09u
mp1 ZN A VDD VDD PMOS_HP L=0.05u W=0.14u
.ENDS 

